CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 110 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
77070354 0
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 943 95 0 1 3
0 2
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9998 0 0
2
43529.9 10
0
2 +V
167 286 312 0 1 3
0 7
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3536 0 0
2
43529.9 9
0
7 Pulser~
4 85 362 0 10 12
0 18 19 8 20 0 0 5 5 5
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4597 0 0
2
43529.9 8
0
9 CC 7-Seg~
183 872 187 0 17 19
10 15 14 13 12 11 10 9 21 2
0 0 0 1 1 1 1 2
0
0 0 21104 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3835 0 0
2
43529.9 7
0
9 2-In AND~
219 677 264 0 3 22
0 16 4 17
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3670 0 0
2
43529.9 6
0
9 2-In AND~
219 509 256 0 3 22
0 6 5 16
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5616 0 0
2
43529.9 5
0
6 74112~
219 749 391 0 7 32
0 7 17 8 17 7 22 3
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
9323 0 0
2
43529.9 4
0
6 74112~
219 602 389 0 7 32
0 7 16 8 16 7 23 4
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
317 0 0
2
43529.9 3
0
6 74112~
219 433 392 0 7 32
0 7 6 8 6 7 24 5
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
3108 0 0
2
43529.9 2
0
6 74112~
219 286 392 0 7 32
0 7 7 8 7 7 25 6
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2A
21 -62 42 -54
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
4299 0 0
2
43529.9 1
0
6 74LS48
188 953 378 0 14 29
0 3 4 5 6 26 27 9 10 11
12 13 14 15 28
0
0 0 4832 0
6 74LS48
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9672 0 0
2
43529.9 0
0
38
6 0 0 0 0 0 0 8 0 0 4 2
632 371
633 371
1 9 2 0 0 0 0 1 4 0 0 4
943 103
943 126
872 126
872 145
0 1 3 0 0 0 0 0 11 8 0 5
790 355
790 490
886 490
886 342
921 342
0 2 4 0 0 16 0 0 11 30 0 5
633 353
633 501
894 501
894 351
921 351
0 3 5 0 0 0 0 0 11 28 0 6
484 356
472 356
472 514
900 514
900 360
921 360
0 4 6 0 0 0 0 0 11 38 0 5
324 356
324 523
907 523
907 369
921 369
0 1 7 0 0 0 0 0 2 25 0 5
230 356
229 356
229 329
286 329
286 321
7 0 3 0 0 0 0 7 0 0 0 2
773 355
803 355
1 0 7 0 0 0 0 2 0 0 13 2
286 321
286 321
0 0 7 0 0 0 0 0 0 13 16 2
347 321
347 419
1 1 7 0 0 0 0 8 7 0 0 4
602 326
602 321
749 321
749 328
1 1 7 0 0 0 0 9 8 0 0 4
433 329
433 321
602 321
602 326
1 1 7 0 0 0 0 10 9 0 0 4
286 329
286 321
433 321
433 329
5 5 7 0 0 0 0 8 7 0 0 4
602 401
602 420
749 420
749 403
5 5 7 0 0 0 0 9 8 0 0 4
433 404
433 420
602 420
602 401
5 5 7 0 0 0 0 10 9 0 0 4
286 404
286 419
433 419
433 404
3 0 8 0 0 0 0 3 0 0 35 4
109 353
132 353
132 454
205 454
7 7 9 0 0 0 0 11 4 0 0 5
985 342
1017 342
1017 286
887 286
887 223
8 6 10 0 0 0 0 11 4 0 0 5
985 351
1012 351
1012 293
881 293
881 223
9 5 11 0 0 0 0 11 4 0 0 5
985 360
1007 360
1007 279
875 279
875 223
10 4 12 0 0 0 0 11 4 0 0 5
985 369
1002 369
1002 272
869 272
869 223
11 3 13 0 0 0 0 11 4 0 0 5
985 378
997 378
997 264
863 264
863 223
12 2 14 0 0 0 0 11 4 0 0 5
985 387
992 387
992 257
857 257
857 223
13 1 15 0 0 0 0 11 4 0 0 5
985 396
987 396
987 249
851 249
851 223
4 2 7 0 0 0 0 10 10 0 0 4
262 374
230 374
230 356
262 356
2 0 16 0 0 0 0 8 0 0 27 2
578 353
540 353
0 4 16 0 0 0 0 0 8 29 0 3
540 256
540 371
578 371
2 7 5 0 0 0 0 6 9 0 0 4
485 265
484 265
484 356
457 356
3 1 16 0 0 0 0 6 5 0 0 3
530 256
653 256
653 255
2 7 4 0 0 0 0 5 8 0 0 4
653 273
644 273
644 353
626 353
2 0 17 0 0 0 0 7 0 0 32 2
725 355
704 355
3 4 17 0 0 0 0 5 7 0 0 4
698 264
704 264
704 373
725 373
3 0 8 0 0 0 0 8 0 0 35 3
572 362
559 362
559 455
3 0 8 0 0 0 0 9 0 0 35 3
403 365
387 365
387 455
3 3 8 0 0 0 0 10 7 0 0 6
256 365
205 365
205 455
694 455
694 364
719 364
1 0 6 0 0 0 0 6 0 0 37 3
485 247
367 247
367 356
4 0 6 0 0 0 0 9 0 0 38 3
409 374
367 374
367 356
7 2 6 0 0 0 0 10 9 0 0 2
310 356
409 356
2
-24 0 0 0 400 0 0 0 255 1 2 1 49
8 Terminal
0 0 0 27
14 29 438 59
29 36 422 58
27 VALEROSO, KENNETH LORVIC M.
-29 0 0 0 400 0 0 0 255 1 2 1 49
8 Terminal
0 0 0 35
118 73 921 110
137 82 901 111
35 BINARY 4-BIT SYNCHRONOUS UP COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
